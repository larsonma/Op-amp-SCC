*******************************************************************
* Filename: Prelab2.cir
* Author: Mitchell Larson <larsonma@msoe.edu>
* Date: May 1, 2018
* Provides:
*	- Signal conditioning circiut that ranges a [0:275]mV signal to
*	- a [0:3200]mV signal using an LM324 opamp.
*******************************************************************


*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM324    1 2 3 4 5
*
c1   11 12 2.887E-12
c2    6  7 30.00E-12
dc    5 53 dy
de   54  5 dy
dlp  90 91 dx
dln  92 90 dx
dp    4  3 dx
egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
fb    7 99 poly(5) vb vc ve vlp vln 0 21.22E6 -1E3 1E3 20E6 -20E6
fpos a 0 vlim 1
w2 3 a vlim sw2
.model sw2 iswitch (ron=1 ion=0 ioff=-1u roff=10meg)
w1 a 0 vlim sw1
.model sw1 iswitch (roff=10meg ioff=0 ion=-1u ron=1)
fneg 0 b vlim -1
w3 4 b vlim sw3
.model sw3 iswitch (ron=1 ion=-1u ioff=0 roff=10meg)
w4 b 0 vlim sw4
.model sw4 iswitch (roff=10meg ioff=-1u ion=0 ron=1)
ga    6  0 11 12 188.5E-6
gcm   0  6 10 99 59.61E-9
iee   3 10 dc 15.09E-6
hlim 90  0 vlim 1K
q1   11  2 13 qx
q2   12  1 14 qx
r2    6  9 100.0E3
rc1   4 11 5.305E3
rc2   4 12 5.305E3
re1  13 10 1.845E3
re2  14 10 1.845E3
ree  10 99 13.25E6
ro1   8  5 50
ro2   7 99 25
rp    3  4 9.082E3
vb    9  0 dc 0
vc    3 53 dc 1.500
ve   54  4 dc 0.822
vlim  7  8 dc 0
vlp  91  0 dc 40
vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=166.7)
.ends


***Circuit Description
***simulation technique: time domain at 1K [0:275]mV

***op-amp power
VCC+ 1 0 DC 5
VCC- 2 0 DC 0

***input voltage
VS 5 0 SIN(137.5m, 137.5m, 1K)

***Design resistances
R1 3 0 1K
R2 3 4 11K

***op-amp***
X1 5 3 1 2 4 lm324

***commands to spice
***simulate two periods
.TRAN 0.0001 2m
.PROBE

.END
